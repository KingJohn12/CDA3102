// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
// CREATED		"Thu Nov 05 11:45:52 2020"

module Four(
	Y
);


output wire	[31:0] Y;

wire	[31:0] Y_ALTERA_SYNTHESIZED;




































assign	Y = Y_ALTERA_SYNTHESIZED;
assign	Y_ALTERA_SYNTHESIZED[0] = 0;
assign	Y_ALTERA_SYNTHESIZED[1] = 0;
assign	Y_ALTERA_SYNTHESIZED[2] = 1;
assign	Y_ALTERA_SYNTHESIZED[3] = 0;
assign	Y_ALTERA_SYNTHESIZED[4] = 0;
assign	Y_ALTERA_SYNTHESIZED[5] = 0;
assign	Y_ALTERA_SYNTHESIZED[6] = 0;
assign	Y_ALTERA_SYNTHESIZED[7] = 0;
assign	Y_ALTERA_SYNTHESIZED[8] = 0;
assign	Y_ALTERA_SYNTHESIZED[9] = 0;
assign	Y_ALTERA_SYNTHESIZED[10] = 0;
assign	Y_ALTERA_SYNTHESIZED[11] = 0;
assign	Y_ALTERA_SYNTHESIZED[12] = 0;
assign	Y_ALTERA_SYNTHESIZED[13] = 0;
assign	Y_ALTERA_SYNTHESIZED[14] = 0;
assign	Y_ALTERA_SYNTHESIZED[15] = 0;
assign	Y_ALTERA_SYNTHESIZED[16] = 0;
assign	Y_ALTERA_SYNTHESIZED[17] = 0;
assign	Y_ALTERA_SYNTHESIZED[18] = 0;
assign	Y_ALTERA_SYNTHESIZED[19] = 0;
assign	Y_ALTERA_SYNTHESIZED[20] = 0;
assign	Y_ALTERA_SYNTHESIZED[21] = 0;
assign	Y_ALTERA_SYNTHESIZED[22] = 0;
assign	Y_ALTERA_SYNTHESIZED[23] = 0;
assign	Y_ALTERA_SYNTHESIZED[24] = 0;
assign	Y_ALTERA_SYNTHESIZED[25] = 0;
assign	Y_ALTERA_SYNTHESIZED[26] = 0;
assign	Y_ALTERA_SYNTHESIZED[27] = 0;
assign	Y_ALTERA_SYNTHESIZED[28] = 0;
assign	Y_ALTERA_SYNTHESIZED[29] = 0;
assign	Y_ALTERA_SYNTHESIZED[30] = 0;
assign	Y_ALTERA_SYNTHESIZED[31] = 0;

endmodule
