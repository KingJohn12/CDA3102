// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
// CREATED		"Thu Nov 05 11:41:11 2020"

module MUX32(
	I0,
	I1,
	I2,
	I3,
	I4,
	I5,
	I6,
	I7,
	I8,
	I9,
	I10,
	I11,
	I12,
	I13,
	I14,
	I15,
	I16,
	I17,
	I18,
	I19,
	I20,
	I21,
	I22,
	I23,
	I24,
	I25,
	I26,
	I27,
	I28,
	I29,
	I30,
	I31,
	S,
	Y
);


input wire	I0;
input wire	I1;
input wire	I2;
input wire	I3;
input wire	I4;
input wire	I5;
input wire	I6;
input wire	I7;
input wire	I8;
input wire	I9;
input wire	I10;
input wire	I11;
input wire	I12;
input wire	I13;
input wire	I14;
input wire	I15;
input wire	I16;
input wire	I17;
input wire	I18;
input wire	I19;
input wire	I20;
input wire	I21;
input wire	I22;
input wire	I23;
input wire	I24;
input wire	I25;
input wire	I26;
input wire	I27;
input wire	I28;
input wire	I29;
input wire	I30;
input wire	I31;
input wire	[4:0] S;
output wire	Y;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;
wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	SYNTHESIZED_WIRE_6;
wire	SYNTHESIZED_WIRE_7;
wire	SYNTHESIZED_WIRE_8;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_13;
wire	SYNTHESIZED_WIRE_14;
wire	SYNTHESIZED_WIRE_15;
wire	SYNTHESIZED_WIRE_16;
wire	SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_25;
wire	SYNTHESIZED_WIRE_26;
wire	SYNTHESIZED_WIRE_27;
wire	SYNTHESIZED_WIRE_28;
wire	SYNTHESIZED_WIRE_29;
wire	SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_31;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_39;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_50;
wire	SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_52;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_61;
wire	SYNTHESIZED_WIRE_62;
wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_67;





Decoder_32	b2v_inst(
	.A(S),
	.Q0(SYNTHESIZED_WIRE_66),
	.Q1(SYNTHESIZED_WIRE_67),
	.Q2(SYNTHESIZED_WIRE_0),
	.Q3(SYNTHESIZED_WIRE_1),
	.Q4(SYNTHESIZED_WIRE_2),
	.Q5(SYNTHESIZED_WIRE_3),
	.Q6(SYNTHESIZED_WIRE_4),
	.Q7(SYNTHESIZED_WIRE_5),
	.Q8(SYNTHESIZED_WIRE_6),
	.Q9(SYNTHESIZED_WIRE_7),
	.Q10(SYNTHESIZED_WIRE_8),
	.Q11(SYNTHESIZED_WIRE_9),
	.Q12(SYNTHESIZED_WIRE_10),
	.Q13(SYNTHESIZED_WIRE_11),
	.Q14(SYNTHESIZED_WIRE_12),
	.Q15(SYNTHESIZED_WIRE_13),
	.Q16(SYNTHESIZED_WIRE_14),
	.Q17(SYNTHESIZED_WIRE_15),
	.Q18(SYNTHESIZED_WIRE_16),
	.Q19(SYNTHESIZED_WIRE_17),
	.Q20(SYNTHESIZED_WIRE_18),
	.Q21(SYNTHESIZED_WIRE_19),
	.Q22(SYNTHESIZED_WIRE_28),
	.Q23(SYNTHESIZED_WIRE_29),
	.Q24(SYNTHESIZED_WIRE_30),
	.Q25(SYNTHESIZED_WIRE_31),
	.Q26(SYNTHESIZED_WIRE_32),
	.Q27(SYNTHESIZED_WIRE_33),
	.Q28(SYNTHESIZED_WIRE_34),
	.Q29(SYNTHESIZED_WIRE_35),
	.Q30(SYNTHESIZED_WIRE_36),
	.Q31(SYNTHESIZED_WIRE_37));

assign	SYNTHESIZED_WIRE_21 = SYNTHESIZED_WIRE_0 & I2;

assign	SYNTHESIZED_WIRE_23 = SYNTHESIZED_WIRE_1 & I3;

assign	SYNTHESIZED_WIRE_25 = SYNTHESIZED_WIRE_2 & I4;

assign	SYNTHESIZED_WIRE_24 = SYNTHESIZED_WIRE_3 & I5;

assign	SYNTHESIZED_WIRE_26 = SYNTHESIZED_WIRE_4 & I6;

assign	SYNTHESIZED_WIRE_27 = SYNTHESIZED_WIRE_5 & I7;

assign	SYNTHESIZED_WIRE_38 = SYNTHESIZED_WIRE_6 & I8;

assign	SYNTHESIZED_WIRE_40 = SYNTHESIZED_WIRE_7 & I9;

assign	SYNTHESIZED_WIRE_39 = SYNTHESIZED_WIRE_8 & I10;

assign	SYNTHESIZED_WIRE_41 = SYNTHESIZED_WIRE_9 & I11;

assign	SYNTHESIZED_WIRE_43 = SYNTHESIZED_WIRE_10 & I12;

assign	SYNTHESIZED_WIRE_42 = SYNTHESIZED_WIRE_11 & I13;

assign	SYNTHESIZED_WIRE_44 = SYNTHESIZED_WIRE_12 & I14;

assign	SYNTHESIZED_WIRE_45 = SYNTHESIZED_WIRE_13 & I15;

assign	SYNTHESIZED_WIRE_46 = SYNTHESIZED_WIRE_14 & I16;

assign	SYNTHESIZED_WIRE_48 = SYNTHESIZED_WIRE_15 & I17;

assign	SYNTHESIZED_WIRE_47 = SYNTHESIZED_WIRE_16 & I18;

assign	SYNTHESIZED_WIRE_49 = SYNTHESIZED_WIRE_17 & I19;

assign	SYNTHESIZED_WIRE_51 = SYNTHESIZED_WIRE_18 & I20;

assign	SYNTHESIZED_WIRE_50 = SYNTHESIZED_WIRE_19 & I21;

assign	SYNTHESIZED_WIRE_62 = SYNTHESIZED_WIRE_20 | SYNTHESIZED_WIRE_21 | SYNTHESIZED_WIRE_22 | SYNTHESIZED_WIRE_23 | SYNTHESIZED_WIRE_24 | SYNTHESIZED_WIRE_25 | SYNTHESIZED_WIRE_26 | SYNTHESIZED_WIRE_27;

assign	SYNTHESIZED_WIRE_52 = SYNTHESIZED_WIRE_28 & I22;

assign	SYNTHESIZED_WIRE_53 = SYNTHESIZED_WIRE_29 & I23;

assign	SYNTHESIZED_WIRE_54 = SYNTHESIZED_WIRE_30 & I24;

assign	SYNTHESIZED_WIRE_56 = SYNTHESIZED_WIRE_31 & I25;

assign	SYNTHESIZED_WIRE_55 = SYNTHESIZED_WIRE_32 & I26;

assign	SYNTHESIZED_WIRE_57 = SYNTHESIZED_WIRE_33 & I27;

assign	SYNTHESIZED_WIRE_59 = SYNTHESIZED_WIRE_34 & I28;

assign	SYNTHESIZED_WIRE_58 = SYNTHESIZED_WIRE_35 & I29;

assign	SYNTHESIZED_WIRE_60 = SYNTHESIZED_WIRE_36 & I30;

assign	SYNTHESIZED_WIRE_61 = SYNTHESIZED_WIRE_37 & I31;

assign	SYNTHESIZED_WIRE_65 = SYNTHESIZED_WIRE_38 | SYNTHESIZED_WIRE_39 | SYNTHESIZED_WIRE_40 | SYNTHESIZED_WIRE_41 | SYNTHESIZED_WIRE_42 | SYNTHESIZED_WIRE_43 | SYNTHESIZED_WIRE_44 | SYNTHESIZED_WIRE_45;

assign	SYNTHESIZED_WIRE_63 = SYNTHESIZED_WIRE_46 | SYNTHESIZED_WIRE_47 | SYNTHESIZED_WIRE_48 | SYNTHESIZED_WIRE_49 | SYNTHESIZED_WIRE_50 | SYNTHESIZED_WIRE_51 | SYNTHESIZED_WIRE_52 | SYNTHESIZED_WIRE_53;

assign	SYNTHESIZED_WIRE_64 = SYNTHESIZED_WIRE_54 | SYNTHESIZED_WIRE_55 | SYNTHESIZED_WIRE_56 | SYNTHESIZED_WIRE_57 | SYNTHESIZED_WIRE_58 | SYNTHESIZED_WIRE_59 | SYNTHESIZED_WIRE_60 | SYNTHESIZED_WIRE_61;

assign	Y = SYNTHESIZED_WIRE_62 | SYNTHESIZED_WIRE_63 | SYNTHESIZED_WIRE_64 | SYNTHESIZED_WIRE_65;

assign	SYNTHESIZED_WIRE_20 = SYNTHESIZED_WIRE_66 & I0;

assign	SYNTHESIZED_WIRE_22 = SYNTHESIZED_WIRE_67 & I1;


endmodule
